& 
Comments: 
VJ-1    = vertically justify proportionally to 2800 
VJ-2    = vertically justify proportionally to 2800; with x2 space between systems
VJ-3    = vertically justify proportionally to 2800; use only inter-system space
VJ-4(#,#,etc. ) = vertically justify to 2800; use only space below designated lines in system
VJ-5(#,#,etc. ) = vertically justify to 2800; use only space below designated lines on page  
  For VJ-4 and VJ-5, if a system or line is designated with a plus sign, it means "add space"
  below this line.  The amount of space (in 10ths of interline distance) is given in 
  square parentheses.  
VEX-# = vertically expand by adding specified distance (10ths of interline) between all lines
MTX(#[x],#[x],etc.)   = move text lines for these line numbers, amount in square parentheses
                          is expressed in 10ths of interline distance.  A positive number
                          moves the text line down.  
MFG(#[x],#[x],etc.)   = move figured harmony for these line numbers, amount in square
                          parentheses is expressed in 10ths of interline distance.  A
                          positive number moves the text line down.  
    


& 
source lib = g:/beethoven/bhl/orch/sym3/outputs/score/pages 
destin lib = g:/beethoven/bhl/orch/sym3/editions/beta-2008/score 
blank page = X 46 575 120 This page is blank 
page id header = X 37 1200C 2950 
page id format = Beethoven Symphony No. 3 in Eb Major, Op. 55 - page ~page     (c) by CCARH 2008
Z MPG-global 
Z 1 Ludwig van Beethoven 
Z 2 Symphony No. 3 in Eb Major, Op. 55 
Z 3             
Z 4 Full Score 
Z 5 300 dots/inch
Z 6 14 dots per staff line
Z 7  

Page    Source          Instructions 
------------------------------------------------------------------- 
001     svp-1 
002     01/01           VJ-6(0,28,56,84,143,177,209,244,291,309,346,361,374)
003     01/02           VJ-6(0,84,167,251,396,528,612,696,784,875) 
004     01/03           VJ-6(0,64,127,191,299,377,509,573,636,704,765) 
005     01/04           VJ-6(0,44,87,131,234,288,338,412,512,556,599,646) 
006     01/05           VJ-6(0,44,87,141,234,288,338,412,512,556,599,646) 
007     01/06           VJ-6(0,46,93,149,246,304,357,475,521,568,617,661) 
008     01/07           VJ-6(0,41,83,124,201,252,299,350,425,457,489,522,553)
009     01/08           VJ-6(0,44,87,131,234,288,338,412,512,556,599,646) 
010     01/09           VJ-6(0,34,81,151,234,288,338,412,512,556,599,646) 
011     01/10           VJ-6(0,46,93,139,246,304,357,475,521,568,617,661) 
012     01/11           VJ-6(0,111,221,332,523,634,745,861,969) 
013     01/12           VJ-6(0,41,83,144,221,262,299,350,425,457,489,522,553)
014     01/13           VJ-6(0,44,87,141,234,288,338,412,512,556,599,646) 
015     01/14           VJ-6(0,41,83,124,201,252,299,350,425,457,489,522,553)
016     01/15           VJ-6(0,46,93,139,256,314,367,475,521,568,617,661) 
017     01/16           VJ-6(0,41,83,124,201,252,299,350,425,457,489,522,553)
018     01/17           VJ-6(0,31,58,62,105,109,126,138,221,234,254,281,314,325,335,346)
019     01/18           VJ-6(0,-1,1,5,22,21,20,26,91,102,106,134,148,144,164,164,159,154)
020     01/19           VJ-6(0,81,161,242,383,481,609,689,770,854) 
021     01/20           VJ-6(0,44,87,131,234,288,338,412,512,556,599,646) 
022     01/21           VJ-6(0,3,-4,1,-7,0,-3,6,10,46,44,39,42,46,30,44,44,60,64)
023     01/22           VJ-6(0,-7,-16,-5,-20,-38,-19,-24,-21,-27,1,-6,-13,-1,-10,-32,-25,-42,-50,-36)
024     01/23           VJ-6(0,87,174,281,387,526,613,700,791,876) 
025     01/24           VJ-6(0,63,126,189,316,393,510,573,635,701,761) 
026     01/25           VJ-6(0,59,119,242,315,388,509,568,627,690,747) 
027     01/26           VJ-6(0,59,119,178,301,374,446,566,625,684,746) 
028     01/27           VJ-6(0,4,1,8,1,-11,-23,4,1,5,4,29,45,56,63,55,67,71,65)
029     01/28           VJ-6(0,5,16,39,53,58,74,79,161,165,181,201,208,235,239,244,259)
030     01/29           VJ-6(0,44,87,131,234,288,338,412,512,556,599,646) 
031     01/30           VJ-6(0,41,83,124,201,252,299,350,425,457,489,522,553)
032     01/31           VJ-6(0,4,-1,6,5,8,6,9,14,56,58,55,62,60,44,57,51,57,67)
033     01/32           VJ-6(0,44,87,131,234,288,338,412,512,556,599,646) 
034     01/33           VJ-6(0,44,87,131,234,288,338,412,512,556,599,646) 
035     01/34           VJ-6(0,104,209,371,496,634,739,843,952) 
036     01/35           VJ-6(0,-8,-14,-11,-21,-23,-40,-19,-26,-17,-11,1,14,58,59,49,72,65,59)
037     01/36           VJ-6(0,81,163,244,387,486,609,690,772,858) 
038     01/37           VJ-6(0,44,87,131,234,288,338,412,512,556,599,646) 
039     01/38           VJ-6(0,44,87,131,234,288,338,412,512,556,599,646) 
040     01/39           VJ-6(0,44,87,131,234,288,338,412,512,556,599,646) 
041     01/40           VJ-6(0,41,83,124,201,252,299,350,425,457,489,522,553)
042     01/41           VJ-6(0,41,83,124,201,252,299,350,425,457,489,522,553)
043     01/42           VJ-6(0,44,87,131,234,288,338,412,512,556,599,646) 
044     01/43           VJ-6(0,31,61,120,201,252,299,350,425,457,489,522,553)
045     01/44           VJ-6(0,64,127,191,319,397,509,573,636,704,765) 
046     01/45           VJ-6(0,41,83,124,201,252,299,350,425,457,489,522,553)
047     01/46           VJ-6(0,41,83,124,201,252,299,350,425,457,489,522,553)
048     01/47           VJ-6(0,44,87,131,234,288,338,412,512,556,599,646) 
049     01/48           VJ-6(0,41,83,124,201,252,299,350,425,447,489,522,553)
050     01/49           VJ-6(0,44,77,131,234,288,338,412,512,556,599,646) 
051     01/50           VJ-6(0,0,1,35,42,26,18,35,36,40,46,59,127,129,149,145,154,166)
052     01/51           VJ-6(0,-14,1,-1,-10,-10,-6,28,46,61,97,89,82,65,56,50,61,64,67)
053     01/52           VJ-6(0,46,91,137,242,299,371,474,519,565,613,656) 
054     01/53           VJ-6(0,-12,-22,-31,-52,-44,-39,-41,-44,-46,-3,-6,-14,-5,-7,-15,-14,-18,-21,-29)
055     01/54           VJ-6(0,41,83,124,201,252,299,350,425,457,489,522,553)
056     01/55           VJ-6(0,41,83,124,201,252,299,350,425,457,489,522,553)
057     01/56           VJ-6(0,87,174,321,407,526,613,700,791,876) 
058     01/57           VJ-6(0,31,63,134,201,252,299,350,425,457,489,522,553)
059     01/58           VJ-6(0,44,87,141,234,288,338,412,512,556,599,646) 
060     01/59           VJ-6(0,44,87,131,234,288,338,412,512,556,599,646) 
061     01/60           VJ-6(0,41,73,124,201,252,299,350,425,457,489,522,553)
062     01/61           VJ-6(0,41,83,124,201,252,299,350,425,457,489,522,553)
